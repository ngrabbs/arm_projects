module top(input  logic        clk, reset,
           output logic [31:0] WriteData, DataAdr,
           output logic        MemWrite,
           output logic [31:0] viewPC,
           output logic [31:0] viewInstr,
           output logic [31:0] viewReadData);

  logic [31:0] PC, Instr, ReadData;

  // instantiate processor and memories
  arm arm(clk, reset, PC, Instr, MemWrite, DataAdr,
          WriteData, ReadData);
  imem imem(PC, Instr);
  dmem dmem(clk, MemWrite, DataAdr, WriteData, ReadData);
  assign viewPC = PC;
  assign viewInstr = Instr;
  assign viewReadData = ReadData;

endmodule