module ex4_19(input  logic [3:0] a,
              output logic p, d);
  always_comb
    case (a)
      4'b0000: {p, d} = 2'b00; // 0
      4'b0001: {p, d} = 2'b00; // 1
      4'b0010: {p, d} = 2'b01; // 2
      4'b0011: {p, d} = 2'b11; // 3
      4'b0100: {p, d} = 2'b00; // 4 
      4'b0101: {p, d} = 2'b01; // 5
      4'b0110: {p, d} = 2'b10; // 6
      4'b0111: {p, d} = 2'b01; // 7
      4'b1000: {p, d} = 2'b00; // 8
      4'b1001: {p, d} = 2'b10; // 9
      4'b1010: {p, d} = 2'b00; // 10
      4'b1011: {p, d} = 2'b01; // 11
      4'b1100: {p, d} = 2'b10; // 12
      4'b1101: {p, d} = 2'b01; // 13
      4'b1110: {p, d} = 2'b00; // 14
      4'b1111: {p, d} = 2'b10; // 15
    endcase
endmodule